magic
tech scmos
timestamp 1717074207
<< nwell >>
rect 3 -4 45 28
<< ntransistor >>
rect 18 -18 20 -13
rect 29 -18 31 -13
<< ptransistor >>
rect 18 2 20 17
rect 29 2 31 17
<< ndiffusion >>
rect 9 -17 12 -13
rect 16 -17 18 -13
rect 9 -18 18 -17
rect 20 -18 29 -13
rect 31 -17 33 -13
rect 37 -17 39 -13
rect 31 -18 39 -17
<< pdiffusion >>
rect 9 15 18 17
rect 9 11 11 15
rect 15 11 18 15
rect 9 7 18 11
rect 9 3 11 7
rect 15 3 18 7
rect 9 2 18 3
rect 20 13 29 17
rect 20 9 22 13
rect 26 9 29 13
rect 20 2 29 9
rect 31 15 39 17
rect 31 11 33 15
rect 37 11 39 15
rect 31 8 39 11
rect 31 4 33 8
rect 37 4 39 8
rect 31 2 39 4
<< ndcontact >>
rect 12 -17 16 -13
rect 33 -17 37 -13
<< pdcontact >>
rect 11 11 15 15
rect 11 3 15 7
rect 22 9 26 13
rect 33 11 37 15
rect 33 4 37 8
<< psubstratepcontact >>
rect 12 -26 16 -22
rect 20 -26 24 -22
rect 28 -26 32 -22
<< nsubstratencontact >>
rect 12 21 16 25
rect 22 21 26 25
rect 33 21 37 25
<< polysilicon >>
rect 18 17 20 19
rect 29 17 31 19
rect 18 -13 20 2
rect 29 -13 31 2
rect 18 -20 20 -18
rect 29 -20 31 -18
<< polycontact >>
rect 13 -9 18 -5
rect 24 -9 29 -5
<< metal1 >>
rect 11 21 12 25
rect 16 21 22 25
rect 26 21 33 25
rect 11 7 15 11
rect 22 13 26 21
rect 22 4 26 9
rect 33 8 37 11
rect 11 1 15 3
rect 33 1 37 4
rect 11 -2 37 1
rect 11 -9 13 -5
rect 22 -9 24 -5
rect 33 -13 37 -2
rect 12 -22 16 -17
rect 33 -18 37 -17
rect 11 -26 12 -22
rect 16 -26 20 -22
rect 24 -26 28 -22
rect 32 -26 37 -22
<< labels >>
rlabel nsubstratencontact 23 22 25 23 1 vdd
rlabel polycontact 14 -7 14 -7 1 A
rlabel polycontact 25 -7 25 -7 1 B
rlabel metal1 35 -7 35 -7 1 out
rlabel metal1 19 -24 19 -24 1 gnd
<< end >>
