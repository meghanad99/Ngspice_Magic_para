** Inverter netlist


* Mosfet

mp1 out in Vdd! Vdd! scmosp w=1u l=0.18u m=1
mn1 out in gnd! gnd! scmosn w=1u l=0.18u m=1

.end

