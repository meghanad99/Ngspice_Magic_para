magic
tech scmos
timestamp 1717076024
<< nwell >>
rect 3 -4 45 28
<< ntransistor >>
rect 18 -18 20 -13
rect 29 -18 31 -13
<< ptransistor >>
rect 18 2 20 17
rect 29 2 31 17
<< ndiffusion >>
rect 9 -18 12 -13
rect 16 -18 18 -13
rect 20 -18 29 -13
rect 31 -18 33 -13
rect 37 -18 39 -13
<< pdiffusion >>
rect 9 15 18 17
rect 9 4 11 15
rect 15 4 18 15
rect 9 2 18 4
rect 20 2 29 17
rect 31 14 39 17
rect 31 4 33 14
rect 37 4 39 14
rect 31 2 39 4
<< ndcontact >>
rect 12 -18 16 -13
rect 33 -18 37 -13
<< pdcontact >>
rect 11 4 15 15
rect 33 4 37 14
<< psubstratepcontact >>
rect 12 -26 16 -22
rect 20 -26 24 -22
rect 28 -26 32 -22
<< nsubstratencontact >>
rect 12 21 16 25
rect 22 21 26 25
rect 33 21 37 25
<< polysilicon >>
rect 18 17 20 19
rect 29 17 31 19
rect 18 -13 20 2
rect 29 -13 31 2
rect 18 -20 20 -18
rect 29 -20 31 -18
<< polycontact >>
rect 13 -5 18 -1
rect 24 -5 29 -1
<< genericcontact >>
rect 23 -17 25 -15
<< metal1 >>
rect 11 21 12 25
rect 16 21 22 25
rect 26 21 33 25
rect 11 15 15 21
rect 11 2 15 4
rect 33 14 37 15
rect 11 -5 13 -1
rect 22 -5 24 -1
rect 33 -8 37 4
rect 12 -11 37 -8
rect 12 -13 16 -11
rect 33 -13 37 -11
rect 22 -22 26 -14
rect 11 -26 12 -22
rect 16 -26 20 -22
rect 24 -26 28 -22
rect 32 -26 37 -22
<< labels >>
rlabel nsubstratencontact 23 22 25 23 1 vdd
rlabel metal1 35 -7 35 -7 1 out
rlabel metal1 19 -24 19 -24 1 gnd
rlabel polycontact 14 -3 14 -3 1 A
rlabel polycontact 26 -3 26 -3 1 B
<< end >>
