magic
tech scmos
timestamp 1717670427
<< nwell >>
rect -31 0 49 32
<< ntransistor >>
rect -20 -20 -18 -16
rect -4 -20 -2 -16
rect 4 -20 6 -16
rect 12 -20 14 -16
rect 20 -20 22 -16
rect 36 -20 38 -16
<< ptransistor >>
rect -20 6 -18 14
rect -4 6 -2 21
rect 4 6 6 21
rect 12 6 14 21
rect 20 6 22 21
rect 36 7 38 15
<< ndiffusion >>
rect -21 -20 -20 -16
rect -18 -20 -17 -16
rect -5 -20 -4 -16
rect -2 -20 4 -16
rect 6 -18 12 -16
rect 6 -20 7 -18
rect 11 -20 12 -18
rect 14 -20 20 -16
rect 22 -20 23 -16
rect 35 -20 36 -16
rect 38 -20 39 -16
<< pdiffusion >>
rect -9 15 -4 21
rect -25 13 -20 14
rect -21 8 -20 13
rect -25 6 -20 8
rect -18 12 -13 14
rect -18 7 -17 12
rect -18 6 -13 7
rect -5 10 -4 15
rect -9 6 -4 10
rect -2 16 4 21
rect -2 11 -1 16
rect 3 11 4 16
rect -2 6 4 11
rect 6 15 12 21
rect 6 10 7 15
rect 11 10 12 15
rect 6 6 12 10
rect 14 16 20 21
rect 14 11 15 16
rect 19 11 20 16
rect 14 6 20 11
rect 22 19 27 21
rect 22 14 23 19
rect 22 6 27 14
rect 31 13 36 15
rect 35 8 36 13
rect 31 7 36 8
rect 38 13 43 15
rect 38 8 39 13
rect 38 7 43 8
<< ndcontact >>
rect -25 -20 -21 -16
rect -17 -20 -13 -16
rect -9 -20 -5 -16
rect 7 -22 11 -18
rect 23 -20 27 -16
rect 31 -20 35 -16
rect 39 -20 43 -16
<< pdcontact >>
rect -25 8 -21 13
rect -17 7 -13 12
rect -9 10 -5 15
rect -1 11 3 16
rect 7 10 11 15
rect 15 11 19 16
rect 23 14 27 19
rect 31 8 35 13
rect 39 8 43 13
<< psubstratepcontact >>
rect -25 -28 -21 -24
rect -9 -28 -5 -24
rect -1 -28 3 -24
rect 15 -28 19 -24
rect 27 -28 31 -24
rect 39 -28 43 -24
<< nsubstratencontact >>
rect -25 25 -21 29
rect -11 25 -7 29
rect 6 25 10 29
rect 14 25 18 29
rect 22 25 26 29
rect 30 25 34 29
<< polysilicon >>
rect -4 21 -2 23
rect 4 21 6 23
rect 12 21 14 23
rect 20 21 22 23
rect -20 14 -18 16
rect 36 15 38 17
rect -20 -16 -18 6
rect -4 -16 -2 6
rect 4 1 6 6
rect 5 -3 6 1
rect 4 -16 6 -3
rect 12 -5 14 6
rect 13 -9 14 -5
rect 12 -16 14 -9
rect 20 -16 22 6
rect 36 -16 38 7
rect -20 -22 -18 -20
rect -4 -22 -2 -20
rect 4 -22 6 -20
rect 12 -22 14 -20
rect 20 -22 22 -20
rect 36 -22 38 -20
<< polycontact >>
rect -24 -9 -20 -5
rect -8 -9 -4 -5
rect 1 -3 5 1
rect 9 -9 13 -5
rect 22 1 26 5
rect 38 -5 42 -1
<< metal1 >>
rect -21 25 -11 29
rect -7 25 6 29
rect 10 25 14 29
rect 18 25 22 29
rect 26 25 30 29
rect 34 25 43 29
rect -25 13 -21 25
rect -1 16 3 25
rect -17 5 -13 7
rect 7 19 27 22
rect 7 15 11 19
rect -9 8 -5 10
rect 39 13 43 25
rect 15 10 19 11
rect 7 8 11 10
rect -9 5 11 8
rect -17 -16 -13 1
rect 16 -12 19 10
rect 31 -8 35 8
rect -9 -15 27 -12
rect -9 -16 -5 -15
rect 23 -16 27 -15
rect -25 -24 -21 -20
rect 31 -16 35 -12
rect 7 -24 11 -22
rect 39 -24 43 -20
rect -21 -28 -9 -24
rect -5 -28 -1 -24
rect 3 -28 15 -24
rect 19 -28 27 -24
rect 31 -28 39 -24
<< m2contact >>
rect -17 1 -13 5
rect -24 -9 -20 -5
rect 1 -3 5 1
rect -8 -9 -4 -5
rect 9 -9 13 -5
rect 22 1 26 5
rect 38 -5 42 -1
rect 31 -12 35 -8
<< metal2 >>
rect -17 5 26 7
rect -13 4 22 5
rect 5 -2 19 1
rect 16 -5 38 -2
rect -20 -9 -8 -5
rect 13 -9 31 -8
rect 9 -12 31 -9
<< labels >>
rlabel metal1 2 27 2 27 5 vdd
rlabel metal1 8 -26 8 -26 1 gnd
rlabel metal2 -11 -7 -11 -7 1 A
rlabel metal2 8 -1 8 -1 1 B
rlabel metal2 -12 5 -12 5 1 A_bar
rlabel metal2 27 -10 27 -10 1 B_bar
<< end >>
