*voltage divider*
r1 in out 1k
r2 out gnd 2k
vin in gnd 1v

.control 
op
print out
.endc
.end

